
interface crc_if(input clk,input  rst_n);



endinterface
