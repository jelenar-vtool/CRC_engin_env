package crc_env_pkg;
    import uvm_pkg::*;
    import crc_pkg::*;


   `include "crc_virtual_sequencer.sv"
   `include "crc_env_cfg.sv"
   //`include "crc_covergroup.sv"  
   `include "crc_virtual_sequence.sv"
   `include "crc_scoreboard.sv"
   `include "crc_env.sv"
	
endpackage 

