
//`include "uvm_pkg.sv"

package crc_test_pkg;

    import uvm_pkg::*;
    import crc_pkg::*;
    import crc_env_pkg::*;
    
    `include "uvm_macros.svh" 
    `include "crc_base_test.sv"
 

endpackage 
