
//`include "uvm_pkg.sv"
`include "uvm_macros.svh" 
`include "apb_pkg.sv"
package apb_test_pkg;

import uvm_pkg::*;
import apb_pkg::*;

// * * * You can include different sequences for specific test bellow * * *

endpackage 

//------------------------------------------------------------------------------------------------------------


