`include "vr_basic_test.sv"

