// * * * Add defines structs enums * * * 





`define IF_ADDR_W 32 //addr width in base_test if
`define IF_DATA_W 32 //data width in base_test if


typedef enum {MASTER1} agent_type_enum1;

