
`include "apb_base_test.sv"
`include "apb_extended_test.sv"
`include "apb_rst_test.sv"
`include "apb_base_sqr_test.sv"
`include "apb_random_test.sv"            
`include "apb_emptread_test.sv"
`include "apb_error_test.sv"
