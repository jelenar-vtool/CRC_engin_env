
//`include "uvm_pkg.sv"
`include "uvm_macros.svh" 
`include "apb_pkg.sv"
package apb_env_pkg;

import uvm_pkg::*;
import apb_pkg::*;

`include "apb_env_cfg.sv"
    `include "vitrual_sequencer.sv"
    `include "vitrual_sequence.sv"
`include "apb_coverage.sv"
`include "apb_scoreboard.sv"

`include "apb_env.sv"

`include "apb_test_list.sv"

endpackage 

//------------------------------------------------------------------------------------------------------------


