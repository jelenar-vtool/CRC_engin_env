
//`include "uvm_pkg.sv"
`include "uvm_macros.svh" 
`include "vr_pkg.sv"
package vr_test_pkg;

import uvm_pkg::*;
import vr_pkg::*;

// * * * You can include different sequences for specific test bellow * * *

endpackage 

